../v1/tinyjambu_control.vhd