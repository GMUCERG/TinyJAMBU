../v1/nlfsr.vhd