../v1/tinyjambu_datapath.vhd